// $Id: $
// File name:   tb_tx.sv
// Created:     12/2/2018
// Author:      Cody Mann
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: This is the test bench for the tx module .
