// $Id: $
// File name:   value_registers.sv
// Created:     11/27/2018
// Author:      Cody Mann
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: This is the block of ahp lite slave module that handles all of the internal registering

module value_registers(

  input wire clk,
  input wire n_rst,
  input wire [3:0] val_loc,
  input wire hwrite_reg,
  input wire [31:0] hwdata,
  input wire [1:0] state,
  input wire [2:0] rx_packet,
  input wire rx_data_ready,
  input wire rx_transfer_active,
  input wire rx_error,
  input wire [6:0] buffer_occupancy,
  input wire [7:0] rx_data,
  input wire tx_transfer_active,
  input wire tx_error,
  output wire d_mode,
  output reg get_rx_data,
  output reg store_tx_data,
  output reg [7:0] tx_data,
  output reg [1:0] tx_packet,
  output reg clear,
  output reg [31:0] hrdata
);

// declaring value location signals 
parameter [3:0] BUFFER4 = 4'd0, 
                 BUFFER3 = 4'd1, 
                 BUFFER2 = 4'd2, 
                 BUFFER1 = 4'd3, 
                 STATUS  = 4'd4, 
                 STATUS_LOWER = 4'd5, 
                 STATUS_UPPER = 4'd6, 
                 ERROR = 4'd7, 
                 ERROR_LOWER = 4'd8,
                 ERROR_UPPER = 4'd9,
                 TX_CONTROL = 4'd10,
                 FLUSH_BUFFER = 4'd11, 
                 BUFFER_OCCUP = 4'd12, 
                 DEFAULT = 4'd13; 

// declaring data types for rx_packet type
parameter [2:0]           OUT = 3'd0, 
						  IN = 3'd1, 
						  DATA0 = 3'd2, 
						  DATA1 = 3'd3, 
						  ACK = 3'd4, 
						  NAK = 3'd5, 
						  STALL = 3'd6; 

// declaring data types for tx_packet
parameter [1:0]          ACK_TX = 2'd0, 
						  NAK_TX = 2'd1, 
						  DATA_TX = 2'd2, 
						  STALL_TX = 2'd3; 

// declaring constants for state input 
parameter [1:0]  IDLE = 2'd0,
                 DATA_TRANSFER = 2'd1, 
                 ERR = 2'd2; 

parameter [4:0] BYTE1 = 5'd0, 
				BYTE2 = 5'd1, 
				BYTE3 = 5'd2, 
				BYTE4 = 5'd3, 
				DATA_IDLE = 5'd6,
				R_BYTE1 = 5'd7, 
				R_BYTE2 = 5'd8, 
				R_BYTE3 = 5'd9, 
				R_BYTE4 = 5'd10; 


// internal signals
reg [15:0] status_reg, status_reg_next, error_reg, error_reg_next;
reg [7:0] tx_control_reg, tx_control_reg_next, flush_buffer_reg_next, flush_buffer_reg;
reg [6:0] buffer_occup_reg;
reg clear_buffer_control, clear_tx_control; 
reg [31:0] rx_data_reg, rx_data_next, hwdata_reg, hwdata_next; 
reg [1:0] buffStateNext, buffState, txStateNext, txState;
reg [4:0] data_state_next, data_state_reg, data_state_prev;

/*D_MODE output logic */
assign d_mode = tx_transfer_active;

/* NEXT STATE LOGIC MODULE CODE */

always_comb
begin: FLUSH_BUFFER_CONTROL_STATE_MACHINE_NEXT_STATE_LOGIC

  buffStateNext = buffState; 

  case(buffState)

  	IDLE: begin 

  		if (flush_buffer_reg != 1'b0) begin 

  			buffStateNext = DATA_TRANSFER; 

  		end 
  		else begin  

  			buffStateNext = IDLE; 

  		end 
  	end 

  	DATA_TRANSFER: begin 

  		if ( flush_buffer_reg == 1'b0) begin 

  			buffStateNext = IDLE; 

  		end 
  		else begin 

  			buffStateNext = DATA_TRANSFER; 

  		end 
  	end 
  endcase 
end

always_comb
begin: TX_CONTROL_STATE_MACHINE_NEXT_STATE_LOGIC

  txStateNext = txState; 

  case(buffState)

  	IDLE: begin 

  		if (tx_control_reg != 1'b0) begin 

  			txStateNext = DATA_TRANSFER; 

  		end 
  		else begin  

  			txStateNext = IDLE; 

  		end 
  	end 

  	DATA_TRANSFER: begin 

  		if ( tx_control_reg == 1'b0) begin 

  			txStateNext = IDLE; 

  		end 
  		else begin 

  			txStateNext = DATA_TRANSFER; 

  		end 
  	end 
  endcase 
end


always_comb
begin: FLUSH_BUFFER_CONTROL_REGISTER_NEXT_STATE_LOGIC

  flush_buffer_reg_next = flush_buffer_reg;

  if ( ( hwrite_reg == 1'b1) & (state == DATA_TRANSFER) & (val_loc== FLUSH_BUFFER) ) begin
    flush_buffer_reg_next = hwdata[7:0];
  end
  else if ( clear_buffer_control == 1'b1) begin
    flush_buffer_reg_next = 8'd0;
  end
end

always_comb
begin: STATUS_REGISTER_NEXT_STATE_LOGIC

  status_reg_next = status_reg;

  if ( (rx_data_ready == 1'b1) & ((rx_packet == DATA0) | (rx_packet == DATA1)) ) begin
    status_reg_next[0] = 1'b1;
  end
  else if ( (status_reg == 1'b1) & (buffer_occupancy == 1'b0) ) begin
    status_reg_next[0] = status_reg[0];
  end
  else begin
    status_reg_next[0] = 1'b0;
  end

  if ( rx_packet == IN) begin
    status_reg_next[1] = 1'b1;
  end
  else if ( (status_reg[1] == 1'b1) & (rx_data_ready == 1'b0) )begin
    status_reg_next[1] = status_reg[1];
  end
  else if ( (status_reg[1] == 1'b1 ) & (rx_data_ready == 1'b1) & (rx_packet != IN) ) begin
    status_reg_next[1] = 1'b0;
  end

  if (rx_packet == OUT) begin
    status_reg_next[2] = 1'b1;
  end
  else if ( ( status_reg[2] == 1'b1 ) & (rx_data_ready == 1'b0) ) begin
    status_reg_next[2] = status_reg[2];
  end
  else if ( (status_reg[2] == 1'b1) & (rx_data_ready == 1'b1) & (rx_packet != OUT) ) begin
    status_reg_next[2] = 1'b0;
  end

  if ( rx_packet == ACK) begin
    status_reg_next[3] = 1'b1;
  end
  else if ( ( status_reg[3] == 1'b1) & (rx_data_ready == 1'b0) ) begin
    status_reg_next[3] = status_reg[3];
  end
  else if ( ( status_reg[3] == 1'b1) & (rx_data_ready == 1'b1) & (rx_packet != ACK) ) begin
    status_reg_next[3] = 1'b0;
  end

  if ( rx_packet == NAK) begin
    status_reg_next[4] = 1'b1;
  end
  else if ( ( status_reg[4] == 1'b1) & (rx_data_ready == 1'b0) ) begin
    status_reg_next[4] = status_reg[4];
  end
  else if ( (status_reg[4] == 1'b1) & (rx_data_ready == 1'b1) & (rx_packet != NAK) ) begin
    status_reg_next[4] = 1'b0;
  end

  if ( rx_transfer_active == 1'b1) begin
    status_reg_next[5] = 1'b1;
  end
  else begin
    status_reg_next[5] = 1'b0;
  end

  if (tx_transfer_active == 1'b1) begin
    status_reg_next[6] = 1'b1;
  end
  else begin
    status_reg_next[6] = 1'b0;
  end
end

always_comb
begin: TX_CONTROL_REGISTER_NEXT_STATE_LOGIC

  tx_control_reg_next = tx_control_reg;

  if ( (hwrite_reg == 1'b1) & (state == DATA_TRANSFER) & (TX_CONTROL) ) begin
    tx_control_reg_next = hwdata[7:0];
  end
  else if (clear_tx_control == 1'b1) begin
    tx_control_reg_next = 8'd0;
  end
end

always_comb
begin: ERROR_REGISTER_NEXT_STATE_LOGIC

  error_reg_next = error_reg;

  if ( rx_error == 1'b1) begin
    error_reg_next[0] = 1'b1;
  end
  else if (rx_transfer_active == 1'b0) begin
    error_reg_next[0] = error_reg[0];
  end
  else begin
    error_reg_next[0] = 1'b0;
  end

  if (tx_error == 1'b1) begin
    error_reg_next[8] = 1'b1;
  end
  else if (tx_transfer_active == 1'b0) begin
    error_reg_next[8] = error_reg[8];
  end
  else begin
    error_reg_next[8] = 1'b0;
  end
end

always_comb 
begin: HWDATA_NEXT_STATE

	hwdata_next = hwdata_reg; 

	if ( (data_state_next != DATA_IDLE) & (data_state_reg == DATA_IDLE)) begin 
		hwdata_next = hwdata;
	end 
end 

always_comb
begin: DATA_BUFFER_STATE_MACHINE_NEXT_STATE_LOGIC


	// assigning arbitrary values to prevent latches
	data_state_next = data_state_reg;
	case(data_state_reg) 

		DATA_IDLE: begin
			if (state == DATA_TRANSFER) begin
				if (val_loc == BUFFER4) begin
					if (hwrite_reg == 1'b1) begin 
						data_state_next = BYTE4;
					end 
					else begin 
						data_state_next = R_BYTE4;
					end 
				end
				if (val_loc== BUFFER2) begin
					if (hwrite_reg == 1'b1) begin 
						data_state_next = BYTE2;
					end 
					else begin 
						data_state_next = R_BYTE2;
					end 
				end
				if (val_loc== BUFFER1) begin
					if (hwrite_reg == 1'b1) begin 
						data_state_next = BYTE1;
					end 
					else begin 
						data_state_next = R_BYTE1;
					end 
				end
				else begin
					data_state_next = DATA_IDLE;
				end
			end
		end 

		//write stattes
		BYTE4: begin 
			data_state_next = BYTE3; 
		end 

		BYTE3: begin 
			data_state_next = BYTE2; 
		end 

		BYTE2: begin 
			data_state_next = BYTE1; 
		end 

		BYTE1: begin 
			data_state_next = DATA_IDLE; 
		end 

		//read stattes
		R_BYTE4: begin 
			data_state_next = R_BYTE3; 
		end 

		R_BYTE3: begin 
			data_state_next = R_BYTE2; 
		end 

		R_BYTE2: begin 
			data_state_next = R_BYTE1; 
		end 

		R_BYTE1: begin 
			data_state_next = DATA_IDLE; 
		end 
	endcase // data_state_reg
end

/*OUTPUT LOGIC BLOCKS */
always_comb
begin: OUTPUT_LOGIC_READING

	// assigning arbitrary values to prevent latches
	hrdata = 32'd0;

	if ( ( hwrite_reg == 1'b0 ) & (state == DATA_TRANSFER) ) begin

		case(val_loc)

			BUFFER4: begin
				hrdata = rx_data_reg;
			end // BUFFER4:

			BUFFER3: begin
				hrdata = {8'd0, rx_data_reg[23:0]};
			end // BUFFER3:

			BUFFER2: begin
				hrdata = {16'd0, rx_data_reg[15:0]};
			end

			BUFFER1: begin
				hrdata = {24'd0, rx_data_reg[7:0]};
			end

			STATUS: begin
				hrdata = {16'd0, status_reg};
			end

			STATUS_LOWER: begin
				hrdata = {24'd0, status_reg[7:0]};
			end

			STATUS_UPPER: begin
				hrdata = {16'd0, status_reg[15:8], 8'd0};
			end

			ERROR: begin
				hrdata = {16'd0, error_reg};
			end

			ERROR_LOWER: begin
				hrdata = {24'd0, error_reg[7:0]};
			end

			ERROR_UPPER: begin
				hrdata = {16'd0, error_reg[15:8], 8'd0};
			end

			BUFFER_OCCUP: begin
				hrdata = {24'd0, buffer_occup_reg};
			end

			TX_CONTROL: begin
				hrdata = {24'd0, tx_control_reg};
			end

			FLUSH_BUFFER: begin
				hrdata = {24'd0, flush_buffer_reg};
			end
		endcase
	end 
end

always_comb
begin: DATA_BUFFER_OUTPUT_LOGIC

	// assigning arbitrary values to prevent latches
	get_rx_data = 'd0;
	store_tx_data = 'd0;
	tx_data = 'd0;
	rx_data_next = rx_data_reg;

	if ((data_state_reg == BYTE1) |
		(data_state_reg == BYTE2) |
		(data_state_reg == BYTE3) |
		(data_state_reg == BYTE4)) begin 
		store_tx_data = 1'b1; 
		tx_data = hwdata_reg[7:0]; 
	end 
	else if ((data_state_reg == R_BYTE1) |
		(data_state_reg == R_BYTE2) |
		(data_state_reg == R_BYTE3) |
		(data_state_reg == R_BYTE4)) begin 
		get_rx_data = 1'b1; 
		rx_data_next = {24'd0, rx_data}; 
	end
end

always_comb
begin: FLUSH_BUFFER_CONTROL_STATE_MACHINE_OUTPUT_LOGIC

  clear_buffer_control = 1'b0; 
  clear = 1'b0; 

  case(buffState)

  	DATA_TRANSFER: begin 

  		clear = 1'b1; 
  		clear_buffer_control = 1'b1; 

  	end 
  endcase // buffState
end

always_comb
begin: TX_CONTROL_STATE_MACHINE_OUTPUT_LOGIC

  clear_tx_control = 1'b0; 
  tx_packet = 1'b0; 

  case(txState)

	DATA_TRANSFER: begin 

		if (tx_transfer_active == 1'b0) begin 

			case(tx_control_reg) 

				8'd1: begin

					if (buffer_occup_reg > 7'd0) begin 

							tx_packet = DATA_TX; 

					end 
				end 

				8'd2: begin 

					tx_packet = ACK_TX; 
				end 

				8'd3: begin 

					tx_packet = NAK_TX; 
				end 

				8'd4: begin 

					tx_packet = STALL_TX; 
				end 
			endcase // tx_control_reg
		end 
	end
  endcase // txState
end

/*REGISTER MODULE CODE */
always_ff @ (posedge clk, negedge n_rst)
begin: REGISTER_LOGIC
	// if reset negation is applied
	if (1'b0 == n_rst ) begin
    	status_reg <= 'd0;
    	error_reg <= 'd0;
    	buffer_occup_reg <= 'd0;
    	tx_control_reg <= 'd0;
    	flush_buffer_reg <= 'd0;
    	rx_data_reg <= 'd0;
	end
	else begin
    	status_reg <= status_reg_next;
	    error_reg <= error_reg_next;
	    buffer_occup_reg <= buffer_occupancy;
	    tx_control_reg <= tx_control_reg_next;
	    flush_buffer_reg <= flush_buffer_reg_next;
	    rx_data_reg <= rx_data_next;
	end
end

always_ff @ (posedge clk, negedge n_rst)
begin: FLUSH_BUFFER_CONTROL_STATE_MACHINE_REGISTER
	// if reset negation is applied
	if (1'b0 == n_rst ) begin

    	buffState <= IDLE;

	end
	else begin

    	buffState <= buffStateNext; 

	end
end

always_ff @ (posedge clk, negedge n_rst)
begin: TX_CONTROL_STATE_MACHINE_REGISTER
	// if reset negation is applied
	if (1'b0 == n_rst ) begin

    	txState <= IDLE;

	end
	else begin

    	txState <= txStateNext; 

	end
end

always_ff @ (posedge clk, negedge n_rst)
begin: DATA_BUFFER_STATE_REGISTER_LOGIC
	// if reset negation is applied
	if (1'b0 == n_rst ) begin
    	data_state_reg <= DATA_IDLE;
	end
	else begin
    	data_state_reg <= data_state_next;
    	data_state_prev <= data_state_reg; 
	end
end

always_ff @ (posedge clk, negedge n_rst)
begin: HWDATA_REGISTER
	// if reset negation is applied
	if (1'b0 == n_rst ) begin
    	hwdata_reg <= 32'd0;
	end
	else begin
    	hwdata_reg <= hwdata_next;
	end
end

endmodule // hwdata register 
